// Copyright 2016 Tudor Timisescu (verificationgentleman.com)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.


typedef enum { OKAY, EXOKAY, SLVERR, DECERR } response_kind_e;



class response extends uvm_sequence_item;
  bit [3:0] id;
  response_kind_e kind;

  function new(string name = get_type_name());
    super.new(name);
  endfunction

  `uvm_object_utils(vgm_axi::response)
endclass
